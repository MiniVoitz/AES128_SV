library verilog;
use verilog.vl_types.all;
entity Rcon_pkg is
end Rcon_pkg;
