library verilog;
use verilog.vl_types.all;
entity InvShiftRows_tb is
end InvShiftRows_tb;
