library verilog;
use verilog.vl_types.all;
entity InvSBox_sv_unit is
end InvSBox_sv_unit;
