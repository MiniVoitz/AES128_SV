library verilog;
use verilog.vl_types.all;
entity MixColumns_tb is
end MixColumns_tb;
