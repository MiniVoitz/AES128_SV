library verilog;
use verilog.vl_types.all;
entity InvSBox_tb is
end InvSBox_tb;
