library verilog;
use verilog.vl_types.all;
entity InvSBox_pkg is
end InvSBox_pkg;
