library verilog;
use verilog.vl_types.all;
entity AES128_tb is
end AES128_tb;
