library verilog;
use verilog.vl_types.all;
entity RoundBlock_tb is
end RoundBlock_tb;
