library verilog;
use verilog.vl_types.all;
entity buffer_tb is
end buffer_tb;
