library verilog;
use verilog.vl_types.all;
entity SBox_pkg2 is
end SBox_pkg2;
