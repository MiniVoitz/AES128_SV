library verilog;
use verilog.vl_types.all;
entity SubBytes_tb is
end SubBytes_tb;
