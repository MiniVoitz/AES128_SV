library verilog;
use verilog.vl_types.all;
entity InvMixColumns_tb is
end InvMixColumns_tb;
