library verilog;
use verilog.vl_types.all;
entity AddRound_Key_tb is
end AddRound_Key_tb;
