library verilog;
use verilog.vl_types.all;
entity LastBlock_tb is
end LastBlock_tb;
