library verilog;
use verilog.vl_types.all;
entity Sbox_sv_unit is
end Sbox_sv_unit;
