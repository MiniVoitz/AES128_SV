library verilog;
use verilog.vl_types.all;
entity mult2to1_tb is
end mult2to1_tb;
