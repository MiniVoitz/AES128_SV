library verilog;
use verilog.vl_types.all;
entity SBox_tb is
end SBox_tb;
