library verilog;
use verilog.vl_types.all;
entity InvSubBytes_tb is
end InvSubBytes_tb;
