library verilog;
use verilog.vl_types.all;
entity KeyExpansion_tb_sv_unit is
end KeyExpansion_tb_sv_unit;
