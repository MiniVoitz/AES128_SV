library verilog;
use verilog.vl_types.all;
entity SBox_pkg is
end SBox_pkg;
